.title KiCad schematic
.model __P20 VDMOS PCHAN
.model __P19 VDMOS PCHAN
.model __P22 VDMOS PCHAN
.model __P21 VDMOS PCHAN
.model __N22 VDMOS NCHAN
.model __N21 VDMOS NCHAN
.model __N20 VDMOS NCHAN
.model __N19 VDMOS NCHAN
.model __N18 VDMOS NCHAN
.model __N17 VDMOS NCHAN
.model __P16 VDMOS PCHAN
.model __P15 VDMOS PCHAN
.model __P18 VDMOS PCHAN
.model __P17 VDMOS PCHAN
.model __N16 VDMOS NCHAN
.model __N15 VDMOS NCHAN
.model __P13 VDMOS PCHAN
.model __P10 VDMOS PCHAN
.model __N10 VDMOS NCHAN
.model __N11 VDMOS NCHAN
.model __P11 VDMOS PCHAN
.model __P12 VDMOS PCHAN
.model __N12 VDMOS NCHAN
.model __N13 VDMOS NCHAN
.model __P25 VDMOS PCHAN
.model __N23 VDMOS NCHAN
.model __N24 VDMOS NCHAN
.model __P23 VDMOS PCHAN
.model __P26 VDMOS PCHAN
.model __N25 VDMOS NCHAN
.model __N26 VDMOS NCHAN
.model __P24 VDMOS PCHAN
.model __P28 VDMOS PCHAN
.model __N27 VDMOS NCHAN
.model __N28 VDMOS NCHAN
.model __P27 VDMOS PCHAN
.model __N31 VDMOS NCHAN
.model __N30 VDMOS NCHAN
.model __P30 VDMOS PCHAN
.model __P31 VDMOS PCHAN
.model __P6 VDMOS PCHAN
.model __N6 VDMOS NCHAN
.model __P1 VDMOS PCHAN
.model __N1 VDMOS NCHAN
.model __P2 VDMOS PCHAN
.model __N2 VDMOS NCHAN
.model __P3 VDMOS PCHAN
.model __P8 VDMOS PCHAN
.model __N8 VDMOS NCHAN
.model __N4 VDMOS NCHAN
.model __N3 VDMOS NCHAN
.model __P4 VDMOS PCHAN
.model __N5 VDMOS NCHAN
.model __P5 VDMOS PCHAN
.model __P29 VDMOS PCHAN
.model __N29 VDMOS NCHAN
.model __N14 VDMOS NCHAN
.model __P14 VDMOS PCHAN
.model __N7 VDMOS NCHAN
.model __N9 VDMOS NCHAN
.model __P9 VDMOS PCHAN
.model __P7 VDMOS PCHAN
MP20 DOUT XORnB1 Net-_P19-D_ __P20
MP19 Net-_P19-D_ XORA1 VDD __P19
MP22 DOUT XORnA1 Net-_P21-D_ __P22
MP21 Net-_P21-D_ NAND01 VDD __P21
MN22 Net-_N21-S_ XORnB1 GND __N22
MN21 DOUT XORnA1 Net-_N21-S_ __N21
MN20 Net-_N19-S_ NAND01 GND __N20
MN19 DOUT XORA1 Net-_N19-S_ __N19
MN18 MIDTEST XORnB0 GND __N18
MN17 XORA1 XORnA0 MIDTEST __N17
MP16 MIDTEST2 NAND0O VDD __P16
MP15 XORA1 XORnB0 MIDTEST2 __P15
MP18 MIDTEST4 DOUT VDD __P18
MP17 XORA1 XORnA0 MIDTEST4 __P17
MN16 MIDTEST3 DOUT GND __N16
MN15 XORA1 NAND0O MIDTEST3 __N15
MP13 NAND01 MONITOR VDD __P13
MP10 NAND0O DOUT VDD __P10
MN10 NAND0O DOUT Net-_N10-S_ __N10
MN11 Net-_N10-S_ MONITOR GND __N11
MP11 NAND0O MONITOR VDD __P11
MP12 NAND01 BUFFERED_DIV2 VDD __P12
MN12 NAND01 BUFFERED_DIV2 Net-_N12-S_ __N12
MN13 Net-_N12-S_ MONITOR GND __N13
MP25 XORnA1 XORA1 VDD __P25
MN23 XORnA1 XORA1 GND __N23
TP4 BUFFERED_DIV2 TP
MN24 XORnA0 NAND0O GND __N24
MP23 XORnA0 NAND0O VDD __P23
MP26 XORnB1 NAND01 VDD __P26
MN25 XORnB1 NAND01 GND __N25
MN26 XORnB0 DOUT GND __N26
MP24 XORnB0 DOUT VDD __P24
MP28 NANDTESTOUT BUFFERED_CLK VDD __P28
TP5 NANDTESTOUT ROON
MN27 NANDTESTOUT BUFFERED_DIV2 Net-_N27-S_ __N27
MN28 Net-_N27-S_ BUFFERED_CLK GND __N28
MP27 NANDTESTOUT BUFFERED_DIV2 VDD __P27
MN31 NORTESTOUT BUFFERED_DIV2 GND __N31
MN30 NORTESTOUT BUFFERED_CLK GND __N30
TP7 NORTESTOUT ROON
MP30 NORTESTOUT BUFFERED_CLK Net-_P30-S_ __P30
MP31 Net-_P30-S_ BUFFERED_DIV2 VDD __P31
MP6 MM2 MM1 VDD __P6
MN6 MM2 MM1 GND __N6
MP1 MM0 MONITOR VDD __P1
MN1 MM0 MONITOR GND __N1
MP2 MM1 MM0 VDD __P2
MN2 MM1 MM0 GND __N2
TP1 GND TP
TP2 VDD TP
MP3 MM6 MM5 VDD __P3
MP8 MM5 MM4 VDD __P8
MN8 MM5 MM4 GND __N8
MN4 MM7 MM6 GND __N4
MN3 MM6 MM5 GND __N3
MP4 MM7 MM6 VDD __P4
MN5 MONITOR MM7 GND __N5
LED1 LEDMR VDD LED
R1 LEDMR MONITOR 1k
MP5 MONITOR MM7 VDD __P5
MP29 BUFFERED_CLK MONITOR VDD __P29
MN29 BUFFERED_CLK MONITOR GND __N29
MN14 BUFFERED_DIV2 DOUT GND __N14
TP6 BUFFERED_CLK ROON
MP14 BUFFERED_DIV2 DOUT VDD __P14
MN7 MM4 MM3 GND __N7
MN9 MM3 MM2 GND __N9
MP9 MM3 MM2 VDD __P9
MP7 MM4 MM3 VDD __P7
.end
