.title KiCad schematic
.model __N5 VDMOS NCHAN
.model __P4 VDMOS PCHAN
.model __N4 VDMOS NCHAN
.model __N3 VDMOS NCHAN
.model __P5 VDMOS PCHAN
.model __P3 VDMOS PCHAN
.model __P1 VDMOS PCHAN
.model __P2 VDMOS PCHAN
.model __N1 VDMOS NCHAN
.model __N2 VDMOS NCHAN
MN5 MONITOR MM1 GND __N5
MP4 MM1 MM2 VDD __P4
MN4 MM1 MM2 GND __N4
MN3 MM2 MM3 GND __N3
MP5 MONITOR MM1 VDD __P5
LED1 Net-_LED1-K_ VDD LED
R1 Net-_LED1-K_ MONITOR 1k
TP3 MM1 TP
MP3 MM2 MM3 VDD __P3
MP1 Net-_N1-D_ MONITOR VDD __P1
MP2 MM3 Net-_N1-D_ VDD __P2
MN1 Net-_N1-D_ MONITOR GND __N1
MN2 MM3 Net-_N1-D_ GND __N2
TP1 GND TP
TP2 VDD TP
.end
