.title KiCad schematic
.model __P1 VDMOS PCHAN
.model __N1 VDMOS NCHAN
.model __P2 VDMOS PCHAN
.model __N2 VDMOS NCHAN
.model __P20 VDMOS PCHAN
.model __P22 VDMOS PCHAN
.model __P21 VDMOS PCHAN
.model __P19 VDMOS PCHAN
.model __N21 VDMOS NCHAN
.model __N22 VDMOS NCHAN
.model __N19 VDMOS NCHAN
.model __N20 VDMOS NCHAN
.model __P25 VDMOS PCHAN
.model __N23 VDMOS NCHAN
.model __P24 VDMOS PCHAN
.model __N26 VDMOS NCHAN
.model __P23 VDMOS PCHAN
.model __N24 VDMOS NCHAN
.model __N25 VDMOS NCHAN
.model __P26 VDMOS PCHAN
.model __N16 VDMOS NCHAN
.model __N15 VDMOS NCHAN
.model __P15 VDMOS PCHAN
.model __P16 VDMOS PCHAN
.model __P17 VDMOS PCHAN
.model __P18 VDMOS PCHAN
.model __N17 VDMOS NCHAN
.model __N18 VDMOS NCHAN
.model __N12 VDMOS NCHAN
.model __N13 VDMOS NCHAN
.model __N29 VDMOS NCHAN
.model __P29 VDMOS PCHAN
.model __P14 VDMOS PCHAN
.model __N14 VDMOS NCHAN
.model __N11 VDMOS NCHAN
.model __P12 VDMOS PCHAN
.model __P10 VDMOS PCHAN
.model __N10 VDMOS NCHAN
.model __P13 VDMOS PCHAN
.model __P11 VDMOS PCHAN
.model __P37 VDMOS PCHAN
.model __N37 VDMOS NCHAN
.model __N30 VDMOS NCHAN
.model __N28 VDMOS NCHAN
.model __P31 VDMOS PCHAN
.model __N31 VDMOS NCHAN
.model __P30 VDMOS PCHAN
.model __P28 VDMOS PCHAN
.model __P27 VDMOS PCHAN
.model __N27 VDMOS NCHAN
.model __N3 VDMOS NCHAN
.model __P3 VDMOS PCHAN
.model __P4 VDMOS PCHAN
.model __N4 VDMOS NCHAN
.model __N5 VDMOS NCHAN
.model __P5 VDMOS PCHAN
.model __N32 VDMOS NCHAN
.model __P32 VDMOS PCHAN
.model __P33 VDMOS PCHAN
.model __N34 VDMOS NCHAN
.model __P34 VDMOS PCHAN
.model __N35 VDMOS NCHAN
.model __N6 VDMOS NCHAN
.model __P6 VDMOS PCHAN
MP1 MONITOR MM2 VDD __P1
MN1 MONITOR MM2 GND __N1
TP12 MONITOR ROON
LED1 LEDMR VDD LED
R1 LEDMR MM2 1k
MP2 NET90OFF MM1 VDD __P2
MN2 NET90OFF MM1 GND __N2
TP13 NET90OFF ROON
MP20 DOUT XORnB1 Net-_P19-D_ __P20
MP22 DOUT XORnA1 Net-_P21-D_ __P22
MP21 Net-_P21-D_ NAND01 VDD __P21
MP19 Net-_P19-D_ XORA1 VDD __P19
MN21 DOUT XORnA1 Net-_N21-S_ __N21
MN22 Net-_N21-S_ XORnB1 GND __N22
MN19 DOUT XORA1 Net-_N19-S_ __N19
MN20 Net-_N19-S_ NAND01 GND __N20
MP25 XORnA1 XORA1 VDD __P25
MN23 XORnA1 XORA1 GND __N23
MP24 XORnB0 DOUT VDD __P24
MN26 XORnB0 DOUT GND __N26
MP23 XORnA0 NAND0O VDD __P23
MN24 XORnA0 NAND0O GND __N24
MN25 XORnB1 NAND01 GND __N25
MP26 XORnB1 NAND01 VDD __P26
MN16 MIDTEST3 DOUT GND __N16
MN15 XORA1 NAND0O MIDTEST3 __N15
MP15 XORA1 XORnB0 MIDTEST2 __P15
MP16 MIDTEST2 NAND0O VDD __P16
MP17 XORA1 XORnA0 MIDTEST4 __P17
MP18 MIDTEST4 DOUT VDD __P18
MN17 XORA1 XORnA0 MIDTEST __N17
MN18 MIDTEST XORnB0 GND __N18
MN12 NAND01 BUFFERED_DIV2 Net-_N12-S_ __N12
MN13 Net-_N12-S_ MONITOR GND __N13
TP6 BUFFERED_CLK ROON
MN29 BUFFERED_CLK MONITOR GND __N29
MP29 BUFFERED_CLK MONITOR VDD __P29
MP14 BUFFERED_DIV2 DOUT VDD __P14
MN14 BUFFERED_DIV2 DOUT GND __N14
TP4 BUFFERED_DIV2 TP
MN11 Net-_N10-S_ MONITOR GND __N11
MP12 NAND01 BUFFERED_DIV2 VDD __P12
MP10 NAND0O DOUT VDD __P10
MN10 NAND0O DOUT Net-_N10-S_ __N10
MP13 NAND01 MONITOR VDD __P13
MP11 NAND0O MONITOR VDD __P11
C3 MM2 GND 1000p
MP37 Net-_N37-D_ BUFFERED_CLK VDD __P37
TP1 GND TP
TP2 VDD TP
MN37 Net-_N37-D_ BUFFERED_CLK GND __N37
MN30 NORTESTOUT NORTESTB GND __N30
MN28 Net-_N27-S_ NANDTESTB GND __N28
MP31 Net-_P30-S_ NORTESTA VDD __P31
MN31 NORTESTOUT NORTESTA GND __N31
TP7 NORTESTOUT ROON
MP30 NORTESTOUT NORTESTB Net-_P30-S_ __P30
MP28 NANDTESTOUT NANDTESTB VDD __P28
MP27 NANDTESTOUT NANDTESTA VDD __P27
MN27 NANDTESTOUT NANDTESTA Net-_N27-S_ __N27
MN3 MM0 MM2 GND __N3
MP3 MM0 MM2 VDD __P3
MP4 MM1 MM0 VDD __P4
MN4 MM1 MM0 GND __N4
MN5 MM2 MM1 GND __N5
TP10 MM1 ROON
MP5 MM2 MM1 VDD __P5
C2 MM1 GND 1000p
MN32 XORTESTOUT XORTESTB XORTESTA __N32
MP32 Net-_P32-D_ XORTESTA VDD __P32
R2 VDD XORTESTOUT 100
MP33 XORTESTOUT XORTESTB Net-_P32-D_ __P33
TP5 NANDTESTOUT ROON
MN34 XORTESTOUT XORTESTA XORTESTB __N34
TP3 XORTESTOUT ROON
TP9 MM2 ROON
TP11 MM0 ROON
C1 MM0 GND 1000p
MP34 NET90OFF Net-_N37-D_ Net-_P34-S_ __P34
R3 TGATE GND 200
TP8 TGATE ROON
MN35 NET90OFF BUFFERED_CLK Net-_N35-S_ __N35
MN6 TGATE BUFFERED_CLK Net-_N35-S_ __N6
R4 VDD TGATE 200
MP6 TGATE Net-_N37-D_ Net-_P34-S_ __P6
.end
