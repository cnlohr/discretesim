.title KiCad schematic
.model __N19 VDMOS NCHAN
.model __N21 VDMOS NCHAN
.model __P23 VDMOS PCHAN
.model __P21 VDMOS PCHAN
.model __P19 VDMOS PCHAN
.model __N23 VDMOS NCHAN
.model __P6 VDMOS PCHAN
.model __N6 VDMOS NCHAN
.model __N12 VDMOS NCHAN
.model __P10 VDMOS PCHAN
.model __N10 VDMOS NCHAN
.model __N8 VDMOS NCHAN
.model __P8 VDMOS PCHAN
.model __P12 VDMOS PCHAN
.model __P2 VDMOS PCHAN
.model __N2 VDMOS NCHAN
.model __N4 VDMOS NCHAN
.model __P4 VDMOS PCHAN
.model __N1 VDMOS NCHAN
.model __P1 VDMOS PCHAN
.model __N20 VDMOS NCHAN
.model __N22 VDMOS NCHAN
.model __N3 VDMOS NCHAN
.model __P20 VDMOS PCHAN
.model __P22 VDMOS PCHAN
.model __P3 VDMOS PCHAN
.model __P25 VDMOS PCHAN
.model __P24 VDMOS PCHAN
.model __P28 VDMOS PCHAN
.model __P27 VDMOS PCHAN
.model __N24 VDMOS NCHAN
.model __N27 VDMOS NCHAN
.model __P7 VDMOS PCHAN
.model __P11 VDMOS PCHAN
.model __P13 VDMOS PCHAN
.model __N5 VDMOS NCHAN
.model __N7 VDMOS NCHAN
.model __N11 VDMOS NCHAN
.model __N13 VDMOS NCHAN
.model __P5 VDMOS PCHAN
.model __N25 VDMOS NCHAN
.model __N28 VDMOS NCHAN
.model __N26 VDMOS NCHAN
.model __P26 VDMOS PCHAN
.model __P16 VDMOS PCHAN
.model __N16 VDMOS NCHAN
.model __P18 VDMOS PCHAN
.model __P17 VDMOS PCHAN
.model __N17 VDMOS NCHAN
.model __N18 VDMOS NCHAN
.model __N14 VDMOS NCHAN
.model __P15 VDMOS PCHAN
.model __P14 VDMOS PCHAN
.model __N15 VDMOS NCHAN
.model __D1 D
.model __N9 VDMOS NCHAN
.model __P9 VDMOS PCHAN
.model __N29 VDMOS NCHAN
.model __N32 VDMOS NCHAN
.model __N33 VDMOS NCHAN
.model __N31 VDMOS NCHAN
.model __N30 VDMOS NCHAN
.model __N34 VDMOS NCHAN
.model __N40 VDMOS NCHAN
.model __N36 VDMOS NCHAN
.model __N38 VDMOS NCHAN
.model __N35 VDMOS NCHAN
.model __N37 VDMOS NCHAN
.model __N39 VDMOS NCHAN
MN19 Net-_N19-D_ nCKO0 GND __N19
MN21 CKMID nFAST Net-_N19-D_ __N21
MP23 nFAST FAST VDD __P23
TP1 nFAST ROON
MP21 Net-_P19-S_ nCKO0 VDD __P21
MP19 CKMID FAST Net-_P19-S_ __P19
MN23 nFAST FAST GND __N23
MP6 Net-_N6-D_ Net-_N4-D_ VDD __P6
MN6 Net-_N6-D_ Net-_N4-D_ GND __N6
MN12 FAST Net-_N10-D_ GND __N12
MP10 Net-_N10-D_ Net-_N10-G_ VDD __P10
MN10 Net-_N10-D_ Net-_N10-G_ GND __N10
MN8 Net-_N10-G_ Net-_N6-D_ GND __N8
MP8 Net-_N10-G_ Net-_N6-D_ VDD __P8
TP5 FAST ROON
MP12 FAST Net-_N10-D_ VDD __P12
C2 GND Net-_N1-D_ 500p
MP2 Net-_N2-D_ Net-_N1-D_ VDD __P2
MN2 Net-_N2-D_ Net-_N1-D_ GND __N2
MN4 Net-_N4-D_ Net-_N2-D_ GND __N4
MP4 Net-_N4-D_ Net-_N2-D_ VDD __P4
MN1 Net-_N1-D_ FAST GND __N1
MP1 Net-_N1-D_ FAST VDD __P1
C1 GND Net-_N2-D_ 500p
MN20 CKO0 FAST Net-_N20-S_ __N20
MN22 Net-_N20-S_ CKMID GND __N22
MN3 nCKO0 CKO0 GND __N3
MP20 Net-_P20-D_ CKMID VDD __P20
MP22 CKO0 nFAST Net-_P20-D_ __P22
MP3 nCKO0 CKO0 VDD __P3
MP25 Net-_N24-D_ CKO2 Net-_P24-D_ __P25
MP24 Net-_P24-D_ nCKO3 VDD __P24
MP28 CKO3 nCKO2 Net-_P27-D_ __P28
MP27 Net-_P27-D_ Net-_N24-D_ VDD __P27
MN24 Net-_N24-D_ nCKO2 Net-_N24-S_ __N24
MN27 CKO3 CKO2 Net-_N27-S_ __N27
MP7 CKO1Mid CKO0 Net-_P5-D_ __P7
MP11 Net-_P11-D_ CKO1Mid VDD __P11
MP13 CKO1 nCKO0 Net-_P11-D_ __P13
MN5 CKO1Mid nCKO0 Net-_N5-S_ __N5
MN7 Net-_N5-S_ nCKO1 GND __N7
MN11 CKO1 CKO0 Net-_N11-S_ __N11
MN13 Net-_N11-S_ CKO1Mid GND __N13
MP5 Net-_P5-D_ nCKO1 VDD __P5
MN25 Net-_N24-S_ nCKO3 GND __N25
MN28 Net-_N27-S_ Net-_N24-D_ GND __N28
MN26 nCKO3 CKO3 GND __N26
MP26 nCKO3 CKO3 VDD __P26
MP16 nCKO2 CKO2 VDD __P16
MN16 nCKO2 CKO2 GND __N16
MP18 CKO2 nCKO1 Net-_P17-D_ __P18
MP17 Net-_P17-D_ Net-_N14-D_ VDD __P17
MN17 CKO2 CKO1 Net-_N17-S_ __N17
MN18 Net-_N17-S_ Net-_N14-D_ GND __N18
MN14 Net-_N14-D_ nCKO1 Net-_N14-S_ __N14
MP15 Net-_N14-D_ CKO1 Net-_P14-D_ __P15
MP14 Net-_P14-D_ nCKO2 VDD __P14
MN15 Net-_N14-S_ nCKO2 GND __N15
D1 Net-_D1-A_ VO __D1
TP3 SW ROON
L2 SW Net-_D1-A_ 4n
MN9 nCKO1 CKO1 GND __N9
MP9 nCKO1 CKO1 VDD __P9
C3 VO GND 1u
TP12 VO ROON
L1 VDD SW 1u
MN29 SW CKO2 GND __N29
TP10 CKO2 ROON
MN32 SW CKO2 GND __N32
MN33 SW CKO2 GND __N33
MN31 SW CKO2 GND __N31
MN30 SW CKO2 GND __N30
MN34 SW CKO2 GND __N34
MN40 SW CKO2 GND __N40
MN36 SW CKO2 GND __N36
MN38 SW CKO2 GND __N38
MN35 SW CKO2 GND __N35
MN37 SW CKO2 GND __N37
MN39 SW CKO2 GND __N39
.end
