.title KiCad schematic
.model __P5 VDMOS PCHAN
.model __P4 VDMOS PCHAN
.model __P6 VDMOS PCHAN
.model __N4 VDMOS NCHAN
.model __N5 VDMOS NCHAN
.model __N6 VDMOS NCHAN
.model __P7 VDMOS PCHAN
.model __N8 VDMOS NCHAN
.model __N7 VDMOS NCHAN
.model __P8 VDMOS PCHAN
.model __D2 D
MP5 MM3 Net-_N4-D_ VDD __P5
MP4 Net-_N4-D_ MONITOR VDD __P4
MP6 MM2 MM3 VDD __P6
MN4 Net-_N4-D_ MONITOR GND __N4
MN5 MM3 Net-_N4-D_ GND __N5
MN6 MM2 MM3 GND __N6
TP_TP2 GND 
TP_TP1 VDD 
R4 Net-_D2-K_ MONITOR 1k
MP7 MM1 MM2 VDD __P7
MN8 MONITOR MM1 GND __N8
TP_TP4 MM1 
MN7 MM1 MM2 GND __N7
MP8 MONITOR MM1 VDD __P8
D2 Net-_D2-K_ VDD __D2
.end
