.title KiCad schematic
.model __P34 VDMOS PCHAN
.model __P6 VDMOS PCHAN
.model __N35 VDMOS NCHAN
.model __N6 VDMOS NCHAN
.model __N37 VDMOS NCHAN
.model __P37 VDMOS PCHAN
.model __N16 VDMOS NCHAN
.model __P15 VDMOS PCHAN
.model __P16 VDMOS PCHAN
.model __N15 VDMOS NCHAN
.model __P1 VDMOS PCHAN
.model __N2 VDMOS NCHAN
.model __P2 VDMOS PCHAN
.model __P7 VDMOS PCHAN
.model __N7 VDMOS NCHAN
.model __P5 VDMOS PCHAN
.model __P4 VDMOS PCHAN
.model __P3 VDMOS PCHAN
.model __N4 VDMOS NCHAN
.model __N3 VDMOS NCHAN
.model __N5 VDMOS NCHAN
.model __N1 VDMOS NCHAN
.model __N29 VDMOS NCHAN
.model __P29 VDMOS PCHAN
.model __P14 VDMOS PCHAN
.model __P13 VDMOS PCHAN
.model __P12 VDMOS PCHAN
.model __N11 VDMOS NCHAN
.model __N14 VDMOS NCHAN
.model __P11 VDMOS PCHAN
.model __N12 VDMOS NCHAN
.model __N13 VDMOS NCHAN
.model __P8 VDMOS PCHAN
.model __P9 VDMOS PCHAN
.model __N10 VDMOS NCHAN
.model __N9 VDMOS NCHAN
.model __N8 VDMOS NCHAN
.model __P10 VDMOS PCHAN
.model __N17 VDMOS NCHAN
.model __N18 VDMOS NCHAN
.model __P17 VDMOS PCHAN
.model __P18 VDMOS PCHAN
MP34 FAST Net-_N37-D_ Net-_P34-S_ __P34
MP6 TGATE Net-_N37-D_ Net-_P34-S_ __P6
MN35 FAST CLK Net-_N35-S_ __N35
MN6 TGATE CLK Net-_N35-S_ __N6
MN37 Net-_N37-D_ CLK GND __N37
TP8 TGATE ROON
R3 TGATE GND 200
MP37 Net-_N37-D_ CLK VDD __P37
R2 VDD TGATE 200
C1 MM0 GND 1000p
C3 MM2 GND 1000p
MN16 Net-_N15-G_ Net-_N16-G_ GND __N16
MP15 Net-_N15-D_ Net-_N15-G_ VDD __P15
MP16 Net-_N15-G_ Net-_N16-G_ VDD __P16
MN15 Net-_N15-D_ Net-_N15-G_ GND __N15
C4 Net-_N15-G_ GND 1000p
R1 LEDMR MM2 1k
MP1 Net-_N1-D_ MM2 VDD __P1
MN2 Net-_N2-D_ MM1 GND __N2
LED1 LEDMR VDD LED
MP2 Net-_N2-D_ MM1 VDD __P2
TP4 CLK90 ROON
MP7 CLK90 Net-_N2-D_ VDD __P7
MN7 CLK90 Net-_N2-D_ GND __N7
C2 MM1 GND 1000p
C5 Net-_N15-D_ GND 1000p
TP11 MM0 ROON
TP9 MM2 ROON
MP5 MM2 MM1 VDD __P5
MP4 MM1 MM0 VDD __P4
MP3 MM0 Net-_N15-D_ VDD __P3
MN4 MM1 MM0 GND __N4
MN3 MM0 Net-_N15-D_ GND __N3
TP10 MM1 ROON
MN5 MM2 MM1 GND __N5
MN1 Net-_N1-D_ MM2 GND __N1
MN29 CLK Net-_N1-D_ GND __N29
MP29 CLK Net-_N1-D_ VDD __P29
TP6 CLK ROON
MP14 Net-_N12-G_ Net-_N11-D_ VDD __P14
MP13 Net-_N13-D_ Net-_N12-D_ VDD __P13
MP12 Net-_N12-D_ Net-_N12-G_ VDD __P12
MN11 Net-_N11-D_ FAST GND __N11
MN14 Net-_N12-G_ Net-_N11-D_ GND __N14
MP11 Net-_N11-D_ FAST VDD __P11
MN12 Net-_N12-D_ Net-_N12-G_ GND __N12
MN13 Net-_N13-D_ Net-_N12-D_ GND __N13
MP8 Net-_N8-D_ Net-_N13-D_ VDD __P8
MP9 Net-_N10-G_ Net-_N8-D_ VDD __P9
MN10 FAST Net-_N10-G_ GND __N10
MN9 Net-_N10-G_ Net-_N8-D_ GND __N9
MN8 Net-_N8-D_ Net-_N13-D_ GND __N8
MP10 FAST Net-_N10-G_ VDD __P10
TP3 FAST ROON
MN17 Net-_N16-G_ Net-_N17-G_ GND __N17
MN18 Net-_N17-G_ MM2 GND __N18
TP2 VDD TP
TP1 GND TP
MP17 Net-_N16-G_ Net-_N17-G_ VDD __P17
MP18 Net-_N17-G_ MM2 VDD __P18
C7 Net-_N17-G_ GND 1000p
C6 Net-_N16-G_ GND 1000p
C8 MM2 GND 1000p
.end
