.title KiCad schematic
.model __P4 VDMOS PCHAN
.model __N5 VDMOS NCHAN
.model __P3 VDMOS PCHAN
.model __P5 VDMOS PCHAN
.model __N3 VDMOS NCHAN
.model __N4 VDMOS NCHAN
.model __P1 VDMOS PCHAN
.model __P2 VDMOS PCHAN
.model __N1 VDMOS NCHAN
.model __N2 VDMOS NCHAN
MP4 MM1 MM2 VDD __P4
MN5 MONITOR MM1 GND __N5
MP3 MM2 MM3 VDD __P3
TP3 MM1 TP
LED1 LEDMR VDD LED
MP5 MONITOR MM1 VDD __P5
R1 LEDMR MONITOR 1k
MN3 MM2 MM3 GND __N3
MN4 MM1 MM2 GND __N4
MP1 MM4 MONITOR VDD __P1
MP2 MM3 MM4 VDD __P2
MN1 MM4 MONITOR GND __N1
MN2 MM3 MM4 GND __N2
TP2 VDD TP
TP1 GND TP
.end
