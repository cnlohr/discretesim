.title KiCad schematic
.model __N25 VDMOS NCHAN
.model __P26 VDMOS PCHAN
.model __P24 VDMOS PCHAN
.model __N26 VDMOS NCHAN
.model __N23 VDMOS NCHAN
.model __P25 VDMOS PCHAN
.model __N24 VDMOS NCHAN
.model __P23 VDMOS PCHAN
.model __N13 VDMOS NCHAN
.model __N12 VDMOS NCHAN
.model __N14 VDMOS NCHAN
.model __P14 VDMOS PCHAN
.model __P19 VDMOS PCHAN
.model __P20 VDMOS PCHAN
.model __N22 VDMOS NCHAN
.model __N21 VDMOS NCHAN
.model __P21 VDMOS PCHAN
.model __P22 VDMOS PCHAN
.model __N20 VDMOS NCHAN
.model __N19 VDMOS NCHAN
.model __N16 VDMOS NCHAN
.model __N15 VDMOS NCHAN
.model __P17 VDMOS PCHAN
.model __P18 VDMOS PCHAN
.model __N18 VDMOS NCHAN
.model __N17 VDMOS NCHAN
.model __P15 VDMOS PCHAN
.model __P16 VDMOS PCHAN
.model __P6 VDMOS PCHAN
.model __P2 VDMOS PCHAN
.model __P1 VDMOS PCHAN
.model __N2 VDMOS NCHAN
.model __N1 VDMOS NCHAN
.model __P3 VDMOS PCHAN
.model __N3 VDMOS NCHAN
.model __P5 VDMOS PCHAN
.model __N5 VDMOS NCHAN
.model __N4 VDMOS NCHAN
.model __P4 VDMOS PCHAN
.model __N6 VDMOS NCHAN
.model __P8 VDMOS PCHAN
.model __P9 VDMOS PCHAN
.model __N9 VDMOS NCHAN
.model __N7 VDMOS NCHAN
.model __N8 VDMOS NCHAN
.model __P7 VDMOS PCHAN
.model __P13 VDMOS PCHAN
.model __P12 VDMOS PCHAN
.model __P10 VDMOS PCHAN
.model __P11 VDMOS PCHAN
.model __N10 VDMOS NCHAN
.model __N11 VDMOS NCHAN
MN25 XORnB1 NAND01 GND __N25
MP26 XORnB1 NAND01 VDD __P26
MP24 XORnB0 XORB0 VDD __P24
MN26 XORnB0 XORB0 GND __N26
MN23 XORnA1 XORA1 GND __N23
MP25 XORnA1 XORA1 VDD __P25
MN24 XORnA0 NAND0O GND __N24
MP23 XORnA0 NAND0O VDD __P23
R3 Net-_N14-D_ NANDA1 1
R2 XORB0 NANDA0 1
MN13 Net-_N12-S_ NANDB1 GND __N13
MN12 NAND01 NANDA1 Net-_N12-S_ __N12
MN14 Net-_N14-D_ XORB0 GND __N14
MP14 Net-_N14-D_ XORB0 VDD __P14
MP19 Net-_P19-D_ XORA1 VDD __P19
MP20 XORB0 XORnB1 Net-_P19-D_ __P20
MN22 Net-_N21-S_ XORnB1 GND __N22
MN21 XORB0 XORnA1 Net-_N21-S_ __N21
MP21 Net-_P21-D_ NAND01 VDD __P21
MP22 XORB0 XORnA1 Net-_P21-D_ __P22
MN20 Net-_N19-S_ NAND01 GND __N20
MN19 XORB0 XORA1 Net-_N19-S_ __N19
R10 XORB0 DOUT 1
MN16 MIDTEST3 XORB0 GND __N16
MN15 XORA1 NAND0O MIDTEST3 __N15
MP17 XORA1 XORnA0 MIDTEST4 __P17
MP18 MIDTEST4 XORB0 VDD __P18
MN18 MIDTEST XORnB0 GND __N18
MN17 XORA1 XORnA0 MIDTEST __N17
MP15 XORA1 XORnB0 MIDTEST2 __P15
MP16 MIDTEST2 NAND0O VDD __P16
MP6 MM2 MM1 VDD __P6
MP2 MM1 MM0 VDD __P2
MP1 MM0 MONITOR VDD __P1
TP1 GND TP
TP2 VDD TP
MN2 MM1 MM0 GND __N2
MN1 MM0 MONITOR GND __N1
MP3 MM6 MM5 VDD __P3
MN3 MM6 MM5 GND __N3
TP3 MM7 TP
MP5 MONITOR MM7 VDD __P5
MN5 MONITOR MM7 GND __N5
MN4 MM7 MM6 GND __N4
MP4 MM7 MM6 VDD __P4
LED1 LEDMR VDD LED
R1 LEDMR MONITOR 1k
MN6 MM2 MM1 GND __N6
MP8 MM5 MM4 VDD __P8
MP9 MM3 MM2 VDD __P9
MN9 MM3 MM2 GND __N9
MN7 MM4 MM3 GND __N7
MN8 MM5 MM4 GND __N8
MP7 MM4 MM3 VDD __P7
R4 MONITOR NANDB0 1
R5 MONITOR NANDB1 1
MP13 NAND01 NANDB1 VDD __P13
MP12 NAND01 NANDA1 VDD __P12
MP10 NAND0O NANDA0 VDD __P10
MP11 NAND0O NANDB0 VDD __P11
MN10 NAND0O NANDA0 Net-_N10-S_ __N10
MN11 Net-_N10-S_ NANDB0 GND __N11
.end
