.title KiCad schematic
.model __P1 VDMOS PCHAN
.model __N1 VDMOS NCHAN
.model __P4 VDMOS PCHAN
.model __P5 VDMOS PCHAN
.model __N4 VDMOS NCHAN
.model __N5 VDMOS NCHAN
.model __P9 VDMOS PCHAN
.model __P10 VDMOS PCHAN
.model __N10 VDMOS NCHAN
.model __N9 VDMOS NCHAN
.model __P8 VDMOS PCHAN
.model __P13 VDMOS PCHAN
.model __N8 VDMOS NCHAN
.model __N13 VDMOS NCHAN
.model __P17 VDMOS PCHAN
.model __N17 VDMOS NCHAN
.model __N18 VDMOS NCHAN
.model __P18 VDMOS PCHAN
.model __N3 VDMOS NCHAN
.model __P3 VDMOS PCHAN
.model __P15 VDMOS PCHAN
.model __N15 VDMOS NCHAN
.model __P16 VDMOS PCHAN
.model __N16 VDMOS NCHAN
.model __N12 VDMOS NCHAN
.model __P12 VDMOS PCHAN
.model __P14 VDMOS PCHAN
.model __P11 VDMOS PCHAN
.model __N14 VDMOS NCHAN
.model __N11 VDMOS NCHAN
.model __N29 VDMOS NCHAN
.model __P29 VDMOS PCHAN
.model __N2 VDMOS NCHAN
.model __P2 VDMOS PCHAN
.model __N7 VDMOS NCHAN
.model __P7 VDMOS PCHAN
.model __N19 VDMOS NCHAN
.model __P19 VDMOS PCHAN
.model __N23 VDMOS NCHAN
.model __N21 VDMOS NCHAN
.model __P6 VDMOS PCHAN
.model __N6 VDMOS NCHAN
.model __P21 VDMOS PCHAN
.model __P23 VDMOS PCHAN
.model __P20 VDMOS PCHAN
.model __P22 VDMOS PCHAN
.model __N22 VDMOS NCHAN
.model __N20 VDMOS NCHAN
C3 MM2 GND 1000p
C5 Net-_N15-D_ GND 1000p
C1 MM0 GND 1000p
MP1 Net-_N1-D_ MM2 VDD __P1
MN1 Net-_N1-D_ MM2 GND __N1
TP9 MM2 ROON
TP11 MM0 ROON
MP4 MM1 MM0 VDD __P4
R1 LEDMR MM2 1k
LED1 LEDMR VDD LED
MP5 MM2 MM1 VDD __P5
MN4 MM1 MM0 GND __N4
MN5 MM2 MM1 GND __N5
TP10 MM1 ROON
MP9 Net-_N10-G_ Net-_N8-D_ VDD __P9
MP10 B Net-_N10-G_ VDD __P10
TP3 B ROON
MN10 B Net-_N10-G_ GND __N10
MN9 Net-_N10-G_ Net-_N8-D_ GND __N9
MP8 Net-_N8-D_ Net-_N13-D_ VDD __P8
MP13 Net-_N13-D_ Net-_N12-D_ VDD __P13
MN8 Net-_N8-D_ Net-_N13-D_ GND __N8
MN13 Net-_N13-D_ Net-_N12-D_ GND __N13
TP1 GND TP
TP2 VDD TP
MP17 Net-_N16-G_ Net-_N17-G_ VDD __P17
MN17 Net-_N16-G_ Net-_N17-G_ GND __N17
C8 MM2 GND 1000p
C7 Net-_N17-G_ GND 1000p
MN18 Net-_N17-G_ MM2 GND __N18
MP18 Net-_N17-G_ MM2 VDD __P18
C6 Net-_N16-G_ GND 1000p
C4 Net-_N15-G_ GND 1000p
MN3 MM0 Net-_N15-D_ GND __N3
MP3 MM0 Net-_N15-D_ VDD __P3
MP15 Net-_N15-D_ Net-_N15-G_ VDD __P15
MN15 Net-_N15-D_ Net-_N15-G_ GND __N15
MP16 Net-_N15-G_ Net-_N16-G_ VDD __P16
MN16 Net-_N15-G_ Net-_N16-G_ GND __N16
MN12 Net-_N12-D_ Net-_N12-G_ GND __N12
MP12 Net-_N12-D_ Net-_N12-G_ VDD __P12
C9 Net-_N12-G_ GND 1000p
MP14 Net-_N12-G_ Net-_N11-D_ VDD __P14
MP11 Net-_N11-D_ B VDD __P11
MN14 Net-_N12-G_ Net-_N11-D_ GND __N14
MN11 Net-_N11-D_ B GND __N11
MN29 A Net-_N1-D_ GND __N29
TP6 A ROON
MP29 A Net-_N1-D_ VDD __P29
MN2 Net-_N2-D_ MM1 GND __N2
MP2 Net-_N2-D_ MM1 VDD __P2
C2 MM1 GND 1000p
MN7 CLK90 Net-_N2-D_ GND __N7
MP7 CLK90 Net-_N2-D_ VDD __P7
TP4 CLK90 ROON
MN19 NB B GND __N19
MP19 NB B VDD __P19
MN23 Net-_N21-D_ NA XOROUT __N23
MN21 Net-_N21-D_ NA B __N21
MP6 NA A VDD __P6
MN6 NA A GND __N6
MP21 XOROUT B Net-_P21-S_ __P21
MP23 A B Net-_P21-S_ __P23
MP20 XOROUT A Net-_P20-S_ __P20
MP22 B A Net-_P20-S_ __P22
TP8 XOROUT ROON
R3 XOROUT GND 200
R2 VDD XOROUT 200
MN22 Net-_N20-D_ A XOROUT __N22
MN20 Net-_N20-D_ A NB __N20
.end
