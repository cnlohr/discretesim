.title KiCad schematic
.model __N1 VDMOS NCHAN
.model __P1 VDMOS PCHAN
.model __N2 VDMOS NCHAN
.model __P2 VDMOS PCHAN
.model __D1 D
.model __N3 VDMOS NCHAN
.model __P3 VDMOS PCHAN
MN1 B0NQ B0S GND __N1
R1 B0NQ B0R 1k
MP1 B0NQ B0S VDD __P1
R2 B0Q B0S 1k
MN2 B0Q B0R GND __N2
MP2 B0Q B0R VDD __P2
D1 B0NQ Net-_D1-A_ __D1
R3 VDD Net-_D1-A_ 1k
MN3 Net-_N3-D_ B0Q GND __N3
MP3 Net-_N3-D_ B0Q VDD __P3
.end
